library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity ROMTriangle367Pts is
		-- Declaro mais um entrada?
		port( noteId : in std_logic_vector(3 downto 0); -- 12 opções - log2(12)= 3.5849625
			  notePt : in std_logic_vector(8 downto 0);
			  DataOut : out std_logic_vector(15 downto 0));
end ROMTriangle367Pts; 

architecture ROM of ROMTriangle367Pts is
	type TROM is array (0 to 15 , 0 to 366) of integer;
		constant value_map : TROM := 
		
-- %%%%%%% MUDO %%%%%%%		
((0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA C3 %%%%%%%	
(-29673, -29346, -29019, -28692, -28365, -28038, -27711, -27384, 
-27057, -26730, -26403, -26076, -25749, -25422, -25095, -24768, 
-24441, -24114, -23787, -23460, -23134, -22807, -22480, -22153, 
-21826, -21499, -21172, -20845, -20518, -20191, -19864, -19537, 
-19210, -18883, -18556, -18229, -17902, -17575, -17248, -16921, 
-16594, -16267, -15940, -15613, -15286, -14959, -14632, -14305, 
-13978, -13651, -13324, -12997, -12670, -12343, -12016, -11689, 
-11362, -11035, -10708, -10381, -10054, -9728, -9401, -9074, 
-8747, -8420, -8093, -7766, -7439, -7112, -6785, -6458, 
-6131, -5804, -5477, -5150, -4823, -4496, -4169, -3842, 
-3515, -3188, -2861, -2534, -2207, -1880, -1553, -1226, 
-899, -572, -245, 82, 409, 736, 1063, 1390, 
1717, 2044, 2371, 2698, 3025, 3351, 3678, 4005, 
4332, 4659, 4986, 5313, 5640, 5967, 6294, 6621, 
6948, 7275, 7602, 7929, 8256, 8583, 8910, 9237, 
9564, 9891, 10218, 10545, 10872, 11199, 11526, 11853, 
12180, 12507, 12834, 13161, 13488, 13815, 14142, 14469, 
14796, 15123, 15450, 15777, 16104, 16431, 16757, 17084, 
17411, 17738, 18065, 18392, 18719, 19046, 19373, 19700, 
20027, 20354, 20681, 21008, 21335, 21662, 21989, 22316, 
22643, 22970, 23297, 23624, 23951, 24278, 24605, 24932, 
25259, 25586, 25913, 26240, 26567, 26894, 27221, 27548, 
27875, 28202, 28529, 28856, 29183, 29510, 29837, 30000, 
29837, 29510, 29183, 28856, 28529, 28202, 27875, 27548, 
27221, 26894, 26567, 26240, 25913, 25586, 25259, 24932, 
24605, 24278, 23951, 23624, 23297, 22970, 22643, 22316, 
21989, 21662, 21335, 21008, 20681, 20354, 20027, 19700, 
19373, 19046, 18719, 18392, 18065, 17738, 17411, 17084, 
16757, 16431, 16104, 15777, 15450, 15123, 14796, 14469, 
14142, 13815, 13488, 13161, 12834, 12507, 12180, 11853, 
11526, 11199, 10872, 10545, 10218, 9891, 9564, 9237, 
8910, 8583, 8256, 7929, 7602, 7275, 6948, 6621, 
6294, 5967, 5640, 5313, 4986, 4659, 4332, 4005, 
3678, 3351, 3025, 2698, 2371, 2044, 1717, 1390, 
1063, 736, 409, 82, -245, -572, -899, -1226, 
-1553, -1880, -2207, -2534, -2861, -3188, -3515, -3842, 
-4169, -4496, -4823, -5150, -5477, -5804, -6131, -6458, 
-6785, -7112, -7439, -7766, -8093, -8420, -8747, -9074, 
-9401, -9728, -10054, -10381, -10708, -11035, -11362, -11689, 
-12016, -12343, -12670, -12997, -13324, -13651, -13978, -14305, 
-14632, -14959, -15286, -15613, -15940, -16267, -16594, -16921, 
-17248, -17575, -17902, -18229, -18556, -18883, -19210, -19537, 
-19864, -20191, -20518, -20845, -21172, -21499, -21826, -22153, 
-22480, -22807, -23134, -23460, -23787, -24114, -24441, -24768, 
-25095, -25422, -25749, -26076, -26403, -26730, -27057, -27384, 
-27711, -28038, -28365, -28692, -29019, -29346, -29673),

-- %%%%%%% NOTA C#3/Db3 %%%%%%%	
(-29653, -29306, -28960, -28613, -28266, -27919, -27572, -27225, 
-26879, -26532, -26185, -25838, -25491, -25145, -24798, -24451, 
-24104, -23757, -23410, -23064, -22717, -22370, -22023, -21676, 
-21329, -20983, -20636, -20289, -19942, -19595, -19249, -18902, 
-18555, -18208, -17861, -17514, -17168, -16821, -16474, -16127, 
-15780, -15434, -15087, -14740, -14393, -14046, -13699, -13353, 
-13006, -12659, -12312, -11965, -11618, -11272, -10925, -10578, 
-10231, -9884, -9538, -9191, -8844, -8497, -8150, -7803, 
-7457, -7110, -6763, -6416, -6069, -5723, -5376, -5029, 
-4682, -4335, -3988, -3642, -3295, -2948, -2601, -2254, 
-1908, -1561, -1214, -867, -520, -173, 173, 520, 
867, 1214, 1561, 1908, 2254, 2601, 2948, 3295, 
3642, 3988, 4335, 4682, 5029, 5376, 5723, 6069, 
6416, 6763, 7110, 7457, 7803, 8150, 8497, 8844, 
9191, 9538, 9884, 10231, 10578, 10925, 11272, 11618, 
11965, 12312, 12659, 13006, 13353, 13699, 14046, 14393, 
14740, 15087, 15434, 15780, 16127, 16474, 16821, 17168, 
17514, 17861, 18208, 18555, 18902, 19249, 19595, 19942, 
20289, 20636, 20983, 21329, 21676, 22023, 22370, 22717, 
23064, 23410, 23757, 24104, 24451, 24798, 25145, 25491, 
25838, 26185, 26532, 26879, 27225, 27572, 27919, 28266, 
28613, 28960, 29306, 29653, 30000, 29653, 29306, 28960, 
28613, 28266, 27919, 27572, 27225, 26879, 26532, 26185, 
25838, 25491, 25145, 24798, 24451, 24104, 23757, 23410, 
23064, 22717, 22370, 22023, 21676, 21329, 20983, 20636, 
20289, 19942, 19595, 19249, 18902, 18555, 18208, 17861, 
17514, 17168, 16821, 16474, 16127, 15780, 15434, 15087, 
14740, 14393, 14046, 13699, 13353, 13006, 12659, 12312, 
11965, 11618, 11272, 10925, 10578, 10231, 9884, 9538, 
9191, 8844, 8497, 8150, 7803, 7457, 7110, 6763, 
6416, 6069, 5723, 5376, 5029, 4682, 4335, 3988, 
3642, 3295, 2948, 2601, 2254, 1908, 1561, 1214, 
867, 520, 173, -173, -520, -867, -1214, -1561, 
-1908, -2254, -2601, -2948, -3295, -3642, -3988, -4335, 
-4682, -5029, -5376, -5723, -6069, -6416, -6763, -7110, 
-7457, -7803, -8150, -8497, -8844, -9191, -9538, -9884, 
-10231, -10578, -10925, -11272, -11618, -11965, -12312, -12659, 
-13006, -13353, -13699, -14046, -14393, -14740, -15087, -15434, 
-15780, -16127, -16474, -16821, -17168, -17514, -17861, -18208, 
-18555, -18902, -19249, -19595, -19942, -20289, -20636, -20983, 
-21329, -21676, -22023, -22370, -22717, -23064, -23410, -23757, 
-24104, -24451, -24798, -25145, -25491, -25838, -26185, -26532, 
-26879, -27225, -27572, -27919, -28266, -28613, -28960, -29306, 
-29653, -30000, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA D3 %%%%%%%	
(-29633, -29266, -28899, -28532, -28165, -27798, -27431, -27064, 
-26697, -26330, -25963, -25596, -25229, -24862, -24495, -24128, 
-23761, -23394, -23028, -22661, -22294, -21927, -21560, -21193, 
-20826, -20459, -20092, -19725, -19358, -18991, -18624, -18257, 
-17890, -17523, -17156, -16789, -16422, -16055, -15688, -15321, 
-14954, -14587, -14220, -13853, -13486, -13119, -12752, -12385, 
-12018, -11651, -11284, -10917, -10550, -10183, -9817, -9450, 
-9083, -8716, -8349, -7982, -7615, -7248, -6881, -6514, 
-6147, -5780, -5413, -5046, -4679, -4312, -3945, -3578, 
-3211, -2844, -2477, -2110, -1743, -1376, -1009, -642, 
-275, 92, 459, 826, 1193, 1560, 1927, 2294, 
2661, 3028, 3394, 3761, 4128, 4495, 4862, 5229, 
5596, 5963, 6330, 6697, 7064, 7431, 7798, 8165, 
8532, 8899, 9266, 9633, 10000, 10367, 10734, 11101, 
11468, 11835, 12202, 12569, 12936, 13303, 13670, 14037, 
14404, 14771, 15138, 15505, 15872, 16239, 16606, 16972, 
17339, 17706, 18073, 18440, 18807, 19174, 19541, 19908, 
20275, 20642, 21009, 21376, 21743, 22110, 22477, 22844, 
23211, 23578, 23945, 24312, 24679, 25046, 25413, 25780, 
26147, 26514, 26881, 27248, 27615, 27982, 28349, 28716, 
29083, 29450, 29817, 30000, 29817, 29450, 29083, 28716, 
28349, 27982, 27615, 27248, 26881, 26514, 26147, 25780, 
25413, 25046, 24679, 24312, 23945, 23578, 23211, 22844, 
22477, 22110, 21743, 21376, 21009, 20642, 20275, 19908, 
19541, 19174, 18807, 18440, 18073, 17706, 17339, 16972, 
16606, 16239, 15872, 15505, 15138, 14771, 14404, 14037, 
13670, 13303, 12936, 12569, 12202, 11835, 11468, 11101, 
10734, 10367, 10000, 9633, 9266, 8899, 8532, 8165, 
7798, 7431, 7064, 6697, 6330, 5963, 5596, 5229, 
4862, 4495, 4128, 3761, 3394, 3028, 2661, 2294, 
1927, 1560, 1193, 826, 459, 92, -275, -642, 
-1009, -1376, -1743, -2110, -2477, -2844, -3211, -3578, 
-3945, -4312, -4679, -5046, -5413, -5780, -6147, -6514, 
-6881, -7248, -7615, -7982, -8349, -8716, -9083, -9450, 
-9817, -10183, -10550, -10917, -11284, -11651, -12018, -12385, 
-12752, -13119, -13486, -13853, -14220, -14587, -14954, -15321, 
-15688, -16055, -16422, -16789, -17156, -17523, -17890, -18257, 
-18624, -18991, -19358, -19725, -20092, -20459, -20826, -21193, 
-21560, -21927, -22294, -22661, -23028, -23394, -23761, -24128, 
-24495, -24862, -25229, -25596, -25963, -26330, -26697, -27064, 
-27431, -27798, -28165, -28532, -28899, -29266, -29633, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA D#3/Eb3 %%%%%%%	
(-29612, -29223, -28835, -28447, -28058, -27670, -27282, -26893, 
-26505, -26117, -25728, -25340, -24951, -24563, -24175, -23786, 
-23398, -23010, -22621, -22233, -21845, -21456, -21068, -20680, 
-20291, -19903, -19515, -19126, -18738, -18350, -17961, -17573, 
-17184, -16796, -16408, -16019, -15631, -15243, -14854, -14466, 
-14078, -13689, -13301, -12913, -12524, -12136, -11748, -11359, 
-10971, -10583, -10194, -9806, -9417, -9029, -8641, -8252, 
-7864, -7476, -7087, -6699, -6311, -5922, -5534, -5146, 
-4757, -4369, -3981, -3592, -3204, -2816, -2427, -2039, 
-1650, -1262, -874, -485, -97, 291, 680, 1068, 
1456, 1845, 2233, 2621, 3010, 3398, 3786, 4175, 
4563, 4951, 5340, 5728, 6117, 6505, 6893, 7282, 
7670, 8058, 8447, 8835, 9223, 9612, 10000, 10388, 
10777, 11165, 11553, 11942, 12330, 12718, 13107, 13495, 
13883, 14272, 14660, 15049, 15437, 15825, 16214, 16602, 
16990, 17379, 17767, 18155, 18544, 18932, 19320, 19709, 
20097, 20485, 20874, 21262, 21650, 22039, 22427, 22816, 
23204, 23592, 23981, 24369, 24757, 25146, 25534, 25922, 
26311, 26699, 27087, 27476, 27864, 28252, 28641, 29029, 
29417, 29806, 30000, 29806, 29417, 29029, 28641, 28252, 
27864, 27476, 27087, 26699, 26311, 25922, 25534, 25146, 
24757, 24369, 23981, 23592, 23204, 22816, 22427, 22039, 
21650, 21262, 20874, 20485, 20097, 19709, 19320, 18932, 
18544, 18155, 17767, 17379, 16990, 16602, 16214, 15825, 
15437, 15049, 14660, 14272, 13883, 13495, 13107, 12718, 
12330, 11942, 11553, 11165, 10777, 10388, 10000, 9612, 
9223, 8835, 8447, 8058, 7670, 7282, 6893, 6505, 
6117, 5728, 5340, 4951, 4563, 4175, 3786, 3398, 
3010, 2621, 2233, 1845, 1456, 1068, 680, 291, 
-97, -485, -874, -1262, -1650, -2039, -2427, -2816, 
-3204, -3592, -3981, -4369, -4757, -5146, -5534, -5922, 
-6311, -6699, -7087, -7476, -7864, -8252, -8641, -9029, 
-9417, -9806, -10194, -10583, -10971, -11359, -11748, -12136, 
-12524, -12913, -13301, -13689, -14078, -14466, -14854, -15243, 
-15631, -16019, -16408, -16796, -17184, -17573, -17961, -18350, 
-18738, -19126, -19515, -19903, -20291, -20680, -21068, -21456, 
-21845, -22233, -22621, -23010, -23398, -23786, -24175, -24563, 
-24951, -25340, -25728, -26117, -26505, -26893, -27282, -27670, 
-28058, -28447, -28835, -29223, -29612, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA E3 %%%%%%%	
(-29588, -29175, -28763, -28351, -27938, -27526, -27113, -26701, 
-26289, -25876, -25464, -25052, -24639, -24227, -23814, -23402, 
-22990, -22577, -22165, -21753, -21340, -20928, -20515, -20103, 
-19691, -19278, -18866, -18454, -18041, -17629, -17216, -16804, 
-16392, -15979, -15567, -15155, -14742, -14330, -13918, -13505, 
-13093, -12680, -12268, -11856, -11443, -11031, -10619, -10206, 
-9794, -9381, -8969, -8557, -8144, -7732, -7320, -6907, 
-6495, -6082, -5670, -5258, -4845, -4433, -4021, -3608, 
-3196, -2784, -2371, -1959, -1546, -1134, -722, -309, 
103, 515, 928, 1340, 1753, 2165, 2577, 2990, 
3402, 3814, 4227, 4639, 5052, 5464, 5876, 6289, 
6701, 7113, 7526, 7938, 8351, 8763, 9175, 9588, 
10000, 10412, 10825, 11237, 11649, 12062, 12474, 12887, 
13299, 13711, 14124, 14536, 14948, 15361, 15773, 16186, 
16598, 17010, 17423, 17835, 18247, 18660, 19072, 19485, 
19897, 20309, 20722, 21134, 21546, 21959, 22371, 22784, 
23196, 23608, 24021, 24433, 24845, 25258, 25670, 26082, 
26495, 26907, 27320, 27732, 28144, 28557, 28969, 29381, 
29794, 30000, 29794, 29381, 28969, 28557, 28144, 27732, 
27320, 26907, 26495, 26082, 25670, 25258, 24845, 24433, 
24021, 23608, 23196, 22784, 22371, 21959, 21546, 21134, 
20722, 20309, 19897, 19485, 19072, 18660, 18247, 17835, 
17423, 17010, 16598, 16186, 15773, 15361, 14948, 14536, 
14124, 13711, 13299, 12887, 12474, 12062, 11649, 11237, 
10825, 10412, 10000, 9588, 9175, 8763, 8351, 7938, 
7526, 7113, 6701, 6289, 5876, 5464, 5052, 4639, 
4227, 3814, 3402, 2990, 2577, 2165, 1753, 1340, 
928, 515, 103, -309, -722, -1134, -1546, -1959, 
-2371, -2784, -3196, -3608, -4021, -4433, -4845, -5258, 
-5670, -6082, -6495, -6907, -7320, -7732, -8144, -8557, 
-8969, -9381, -9794, -10206, -10619, -11031, -11443, -11856, 
-12268, -12680, -13093, -13505, -13918, -14330, -14742, -15155, 
-15567, -15979, -16392, -16804, -17216, -17629, -18041, -18454, 
-18866, -19278, -19691, -20103, -20515, -20928, -21340, -21753, 
-22165, -22577, -22990, -23402, -23814, -24227, -24639, -25052, 
-25464, -25876, -26289, -26701, -27113, -27526, -27938, -28351, 
-28763, -29175, -29588, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA F3 %%%%%%%	
(-29564, -29127, -28691, -28255, -27818, -27382, -26945, -26509, 
-26073, -25636, -25200, -24764, -24327, -23891, -23455, -23018, 
-22582, -22145, -21709, -21273, -20836, -20400, -19964, -19527, 
-19091, -18655, -18218, -17782, -17345, -16909, -16473, -16036, 
-15600, -15164, -14727, -14291, -13855, -13418, -12982, -12545, 
-12109, -11673, -11236, -10800, -10364, -9927, -9491, -9055, 
-8618, -8182, -7745, -7309, -6873, -6436, -6000, -5564, 
-5127, -4691, -4255, -3818, -3382, -2945, -2509, -2073, 
-1636, -1200, -764, -327, 109, 545, 982, 1418, 
1855, 2291, 2727, 3164, 3600, 4036, 4473, 4909, 
5345, 5782, 6218, 6655, 7091, 7527, 7964, 8400, 
8836, 9273, 9709, 10145, 10582, 11018, 11455, 11891, 
12327, 12764, 13200, 13636, 14073, 14509, 14945, 15382, 
15818, 16255, 16691, 17127, 17564, 18000, 18436, 18873, 
19309, 19745, 20182, 20618, 21055, 21491, 21927, 22364, 
22800, 23236, 23673, 24109, 24545, 24982, 25418, 25855, 
26291, 26727, 27164, 27600, 28036, 28473, 28909, 29345, 
29782, 30000, 29782, 29345, 28909, 28473, 28036, 27600, 
27164, 26727, 26291, 25855, 25418, 24982, 24545, 24109, 
23673, 23236, 22800, 22364, 21927, 21491, 21055, 20618, 
20182, 19745, 19309, 18873, 18436, 18000, 17564, 17127, 
16691, 16255, 15818, 15382, 14945, 14509, 14073, 13636, 
13200, 12764, 12327, 11891, 11455, 11018, 10582, 10145, 
9709, 9273, 8836, 8400, 7964, 7527, 7091, 6655, 
6218, 5782, 5345, 4909, 4473, 4036, 3600, 3164, 
2727, 2291, 1855, 1418, 982, 545, 109, -327, 
-764, -1200, -1636, -2073, -2509, -2945, -3382, -3818, 
-4255, -4691, -5127, -5564, -6000, -6436, -6873, -7309, 
-7745, -8182, -8618, -9055, -9491, -9927, -10364, -10800, 
-11236, -11673, -12109, -12545, -12982, -13418, -13855, -14291, 
-14727, -15164, -15600, -16036, -16473, -16909, -17345, -17782, 
-18218, -18655, -19091, -19527, -19964, -20400, -20836, -21273, 
-21709, -22145, -22582, -23018, -23455, -23891, -24327, -24764, 
-25200, -25636, -26073, -26509, -26945, -27382, -27818, -28255, 
-28691, -29127, -29564, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA F#3/Gb3 %%%%%%%	
(-29537, -29073, -28610, -28147, -27683, -27220, -26757, -26293, 
-25830, -25367, -24903, -24440, -23977, -23514, -23050, -22587, 
-22124, -21660, -21197, -20734, -20270, -19807, -19344, -18880, 
-18417, -17954, -17490, -17027, -16564, -16100, -15637, -15174, 
-14710, -14247, -13784, -13320, -12857, -12394, -11931, -11467, 
-11004, -10541, -10077, -9614, -9151, -8687, -8224, -7761, 
-7297, -6834, -6371, -5907, -5444, -4981, -4517, -4054, 
-3591, -3127, -2664, -2201, -1737, -1274, -811, -347, 
116, 579, 1042, 1506, 1969, 2432, 2896, 3359, 
3822, 4286, 4749, 5212, 5676, 6139, 6602, 7066, 
7529, 7992, 8456, 8919, 9382, 9846, 10309, 10772, 
11236, 11699, 12162, 12625, 13089, 13552, 14015, 14479, 
14942, 15405, 15869, 16332, 16795, 17259, 17722, 18185, 
18649, 19112, 19575, 20039, 20502, 20965, 21429, 21892, 
22355, 22819, 23282, 23745, 24208, 24672, 25135, 25598, 
26062, 26525, 26988, 27452, 27915, 28378, 28842, 29305, 
29768, 30000, 29768, 29305, 28842, 28378, 27915, 27452, 
26988, 26525, 26062, 25598, 25135, 24672, 24208, 23745, 
23282, 22819, 22355, 21892, 21429, 20965, 20502, 20039, 
19575, 19112, 18649, 18185, 17722, 17259, 16795, 16332, 
15869, 15405, 14942, 14479, 14015, 13552, 13089, 12625, 
12162, 11699, 11236, 10772, 10309, 9846, 9382, 8919, 
8456, 7992, 7529, 7066, 6602, 6139, 5676, 5212, 
4749, 4286, 3822, 3359, 2896, 2432, 1969, 1506, 
1042, 579, 116, -347, -811, -1274, -1737, -2201, 
-2664, -3127, -3591, -4054, -4517, -4981, -5444, -5907, 
-6371, -6834, -7297, -7761, -8224, -8687, -9151, -9614, 
-10077, -10541, -11004, -11467, -11931, -12394, -12857, -13320, 
-13784, -14247, -14710, -15174, -15637, -16100, -16564, -17027, 
-17490, -17954, -18417, -18880, -19344, -19807, -20270, -20734, 
-21197, -21660, -22124, -22587, -23050, -23514, -23977, -24440, 
-24903, -25367, -25830, -26293, -26757, -27220, -27683, -28147, 
-28610, -29073, -29537, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA G3 %%%%%%%	
(-29510, -29020, -28531, -28041, -27551, -27061, -26571, -26082, 
-25592, -25102, -24612, -24122, -23633, -23143, -22653, -22163, 
-21673, -21184, -20694, -20204, -19714, -19224, -18735, -18245, 
-17755, -17265, -16776, -16286, -15796, -15306, -14816, -14327, 
-13837, -13347, -12857, -12367, -11878, -11388, -10898, -10408, 
-9918, -9429, -8939, -8449, -7959, -7469, -6980, -6490, 
-6000, -5510, -5020, -4531, -4041, -3551, -3061, -2571, 
-2082, -1592, -1102, -612, -122, 367, 857, 1347, 
1837, 2327, 2816, 3306, 3796, 4286, 4776, 5265, 
5755, 6245, 6735, 7224, 7714, 8204, 8694, 9184, 
9673, 10163, 10653, 11143, 11633, 12122, 12612, 13102, 
13592, 14082, 14571, 15061, 15551, 16041, 16531, 17020, 
17510, 18000, 18490, 18980, 19469, 19959, 20449, 20939, 
21429, 21918, 22408, 22898, 23388, 23878, 24367, 24857, 
25347, 25837, 26327, 26816, 27306, 27796, 28286, 28776, 
29265, 29755, 30000, 29755, 29265, 28776, 28286, 27796, 
27306, 26816, 26327, 25837, 25347, 24857, 24367, 23878, 
23388, 22898, 22408, 21918, 21429, 20939, 20449, 19959, 
19469, 18980, 18490, 18000, 17510, 17020, 16531, 16041, 
15551, 15061, 14571, 14082, 13592, 13102, 12612, 12122, 
11633, 11143, 10653, 10163, 9673, 9184, 8694, 8204, 
7714, 7224, 6735, 6245, 5755, 5265, 4776, 4286, 
3796, 3306, 2816, 2327, 1837, 1347, 857, 367, 
-122, -612, -1102, -1592, -2082, -2571, -3061, -3551, 
-4041, -4531, -5020, -5510, -6000, -6490, -6980, -7469, 
-7959, -8449, -8939, -9429, -9918, -10408, -10898, -11388, 
-11878, -12367, -12857, -13347, -13837, -14327, -14816, -15306, 
-15796, -16286, -16776, -17265, -17755, -18245, -18735, -19224, 
-19714, -20204, -20694, -21184, -21673, -22163, -22653, -23143, 
-23633, -24122, -24612, -25102, -25592, -26082, -26571, -27061, 
-27551, -28041, -28531, -29020, -29510, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA G#3/Ab3 %%%%%%%	
(-29481, -28961, -28442, -27922, -27403, -26883, -26364, -25844, 
-25325, -24805, -24286, -23766, -23247, -22727, -22208, -21688, 
-21169, -20649, -20130, -19610, -19091, -18571, -18052, -17532, 
-17013, -16494, -15974, -15455, -14935, -14416, -13896, -13377, 
-12857, -12338, -11818, -11299, -10779, -10260, -9740, -9221, 
-8701, -8182, -7662, -7143, -6623, -6104, -5584, -5065, 
-4545, -4026, -3506, -2987, -2468, -1948, -1429, -909, 
-390, 130, 649, 1169, 1688, 2208, 2727, 3247, 
3766, 4286, 4805, 5325, 5844, 6364, 6883, 7403, 
7922, 8442, 8961, 9481, 10000, 10519, 11039, 11558, 
12078, 12597, 13117, 13636, 14156, 14675, 15195, 15714, 
16234, 16753, 17273, 17792, 18312, 18831, 19351, 19870, 
20390, 20909, 21429, 21948, 22468, 22987, 23506, 24026, 
24545, 25065, 25584, 26104, 26623, 27143, 27662, 28182, 
28701, 29221, 29740, 30000, 29740, 29221, 28701, 28182, 
27662, 27143, 26623, 26104, 25584, 25065, 24545, 24026, 
23506, 22987, 22468, 21948, 21429, 20909, 20390, 19870, 
19351, 18831, 18312, 17792, 17273, 16753, 16234, 15714, 
15195, 14675, 14156, 13636, 13117, 12597, 12078, 11558, 
11039, 10519, 10000, 9481, 8961, 8442, 7922, 7403, 
6883, 6364, 5844, 5325, 4805, 4286, 3766, 3247, 
2727, 2208, 1688, 1169, 649, 130, -390, -909, 
-1429, -1948, -2468, -2987, -3506, -4026, -4545, -5065, 
-5584, -6104, -6623, -7143, -7662, -8182, -8701, -9221, 
-9740, -10260, -10779, -11299, -11818, -12338, -12857, -13377, 
-13896, -14416, -14935, -15455, -15974, -16494, -17013, -17532, 
-18052, -18571, -19091, -19610, -20130, -20649, -21169, -21688, 
-22208, -22727, -23247, -23766, -24286, -24805, -25325, -25844, 
-26364, -26883, -27403, -27922, -28442, -28961, -29481, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA A3 %%%%%%%	
(-29450, -28899, -28349, -27798, -27248, -26697, -26147, -25596, 
-25046, -24495, -23945, -23394, -22844, -22294, -21743, -21193, 
-20642, -20092, -19541, -18991, -18440, -17890, -17339, -16789, 
-16239, -15688, -15138, -14587, -14037, -13486, -12936, -12385, 
-11835, -11284, -10734, -10183, -9633, -9083, -8532, -7982, 
-7431, -6881, -6330, -5780, -5229, -4679, -4128, -3578, 
-3028, -2477, -1927, -1376, -826, -275, 275, 826, 
1376, 1927, 2477, 3028, 3578, 4128, 4679, 5229, 
5780, 6330, 6881, 7431, 7982, 8532, 9083, 9633, 
10183, 10734, 11284, 11835, 12385, 12936, 13486, 14037, 
14587, 15138, 15688, 16239, 16789, 17339, 17890, 18440, 
18991, 19541, 20092, 20642, 21193, 21743, 22294, 22844, 
23394, 23945, 24495, 25046, 25596, 26147, 26697, 27248, 
27798, 28349, 28899, 29450, 30000, 29450, 28899, 28349, 
27798, 27248, 26697, 26147, 25596, 25046, 24495, 23945, 
23394, 22844, 22294, 21743, 21193, 20642, 20092, 19541, 
18991, 18440, 17890, 17339, 16789, 16239, 15688, 15138, 
14587, 14037, 13486, 12936, 12385, 11835, 11284, 10734, 
10183, 9633, 9083, 8532, 7982, 7431, 6881, 6330, 
5780, 5229, 4679, 4128, 3578, 3028, 2477, 1927, 
1376, 826, 275, -275, -826, -1376, -1927, -2477, 
-3028, -3578, -4128, -4679, -5229, -5780, -6330, -6881, 
-7431, -7982, -8532, -9083, -9633, -10183, -10734, -11284, 
-11835, -12385, -12936, -13486, -14037, -14587, -15138, -15688, 
-16239, -16789, -17339, -17890, -18440, -18991, -19541, -20092, 
-20642, -21193, -21743, -22294, -22844, -23394, -23945, -24495, 
-25046, -25596, -26147, -26697, -27248, -27798, -28349, -28899, 
-29450, -30000, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA A#3/Bb3 %%%%%%%	
(-29417, -28835, -28252, -27670, -27087, -26505, -25922, -25340, 
-24757, -24175, -23592, -23010, -22427, -21845, -21262, -20680, 
-20097, -19515, -18932, -18350, -17767, -17184, -16602, -16019, 
-15437, -14854, -14272, -13689, -13107, -12524, -11942, -11359, 
-10777, -10194, -9612, -9029, -8447, -7864, -7282, -6699, 
-6117, -5534, -4951, -4369, -3786, -3204, -2621, -2039, 
-1456, -874, -291, 291, 874, 1456, 2039, 2621, 
3204, 3786, 4369, 4951, 5534, 6117, 6699, 7282, 
7864, 8447, 9029, 9612, 10194, 10777, 11359, 11942, 
12524, 13107, 13689, 14272, 14854, 15437, 16019, 16602, 
17184, 17767, 18350, 18932, 19515, 20097, 20680, 21262, 
21845, 22427, 23010, 23592, 24175, 24757, 25340, 25922, 
26505, 27087, 27670, 28252, 28835, 29417, 30000, 29417, 
28835, 28252, 27670, 27087, 26505, 25922, 25340, 24757, 
24175, 23592, 23010, 22427, 21845, 21262, 20680, 20097, 
19515, 18932, 18350, 17767, 17184, 16602, 16019, 15437, 
14854, 14272, 13689, 13107, 12524, 11942, 11359, 10777, 
10194, 9612, 9029, 8447, 7864, 7282, 6699, 6117, 
5534, 4951, 4369, 3786, 3204, 2621, 2039, 1456, 
874, 291, -291, -874, -1456, -2039, -2621, -3204, 
-3786, -4369, -4951, -5534, -6117, -6699, -7282, -7864, 
-8447, -9029, -9612, -10194, -10777, -11359, -11942, -12524, 
-13107, -13689, -14272, -14854, -15437, -16019, -16602, -17184, 
-17767, -18350, -18932, -19515, -20097, -20680, -21262, -21845, 
-22427, -23010, -23592, -24175, -24757, -25340, -25922, -26505, 
-27087, -27670, -28252, -28835, -29417, -30000, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- %%%%%%% NOTA B3 %%%%%%%	
(-29381, -28763, -28144, -27526, -26907, -26289, -25670, -25052, 
-24433, -23814, -23196, -22577, -21959, -21340, -20722, -20103, 
-19485, -18866, -18247, -17629, -17010, -16392, -15773, -15155, 
-14536, -13918, -13299, -12680, -12062, -11443, -10825, -10206, 
-9588, -8969, -8351, -7732, -7113, -6495, -5876, -5258, 
-4639, -4021, -3402, -2784, -2165, -1546, -928, -309, 
309, 928, 1546, 2165, 2784, 3402, 4021, 4639, 
5258, 5876, 6495, 7113, 7732, 8351, 8969, 9588, 
10206, 10825, 11443, 12062, 12680, 13299, 13918, 14536, 
15155, 15773, 16392, 17010, 17629, 18247, 18866, 19485, 
20103, 20722, 21340, 21959, 22577, 23196, 23814, 24433, 
25052, 25670, 26289, 26907, 27526, 28144, 28763, 29381, 
30000, 29381, 28763, 28144, 27526, 26907, 26289, 25670, 
25052, 24433, 23814, 23196, 22577, 21959, 21340, 20722, 
20103, 19485, 18866, 18247, 17629, 17010, 16392, 15773, 
15155, 14536, 13918, 13299, 12680, 12062, 11443, 10825, 
10206, 9588, 8969, 8351, 7732, 7113, 6495, 5876, 
5258, 4639, 4021, 3402, 2784, 2165, 1546, 928, 
309, -309, -928, -1546, -2165, -2784, -3402, -4021, 
-4639, -5258, -5876, -6495, -7113, -7732, -8351, -8969, 
-9588, -10206, -10825, -11443, -12062, -12680, -13299, -13918, 
-14536, -15155, -15773, -16392, -17010, -17629, -18247, -18866, 
-19485, -20103, -20722, -21340, -21959, -22577, -23196, -23814, 
-24433, -25052, -25670, -26289, -26907, -27526, -28144, -28763, 
-29381, -30000, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

-- DE MODO A ENCHER O ARRAY PARA BASE 2
(0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

(0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0),

(0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0));

		
	begin
		DataOut <= std_logic_vector(to_signed(value_map(to_integer(unsigned(noteId)), to_integer(unsigned(notePt))), 16));
end ROM;